`timescale 1ns / 1ps

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
   // ��Ƽ�÷��� 2�� �ް� 1�� ��� 2x1
   
   module mux_2_1(
            input [1:0] d,
            input s,
            output f);
            
            assign f =s ? d[1] :d[0];
            
   endmodule  
   
   
      ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
   // ��Ƽ�÷���4x1
   
   module mux_4_1(
            input [3:0] d,
            input [1:0] s, //s�� ���� ���� ��µǴ� d�� ��Ʈ�� �޶���
            output f);
            
            assign f = d[s];
            
   endmodule  
   
         ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
   // ��Ƽ�÷���8x1
   
   module mux_8_1(
            input [7:0] d,
            input [2:0] s, //s�� ���� ���� ��µǴ� d�� ��Ʈ�� �޶���
            output f);
            
            assign f = d[s];
            
   endmodule  
   
 ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
   // ���Ƽ�÷���1x4
   
   module demux_1_4(
            input d,
            input [1:0] s,
            output [3:0] f);
            
            assign f = (s==2'b00) ? {3'd000, d} : 
                             ((s==2'b01) ? {2'b00, d, 1'b0} :
                             ((s==2'b10) ? {1'b0, d, 2'b00} :{d,3'b000}));
                                                
   endmodule
   
   
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
   // ��Ƽ�÷��� +���Ƽ�÷��� (��Ƽ�÷���)
   
   module mux_demux_test(
                input [3:0] d,
                input [1:0] mux_s, demux_s,
                output [3:0] f);
              
              wire line;
              
              mux_4_1 mux(.d(d), .s(mux_s), .f(line));
              demux_1_4 demux(.d(line), .s(demux_s), .f(f));
  
  endmodule
